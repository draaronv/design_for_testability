library ieee;use ieee.std_logic_1164.all;Entity TriStateBuffer16 is  Port(Data : in std_logic_vector(15 downto 0);       En : in std_logic;       Outp : out std_logic_vector(15 downto 0));end;Architecture behav of TriStateBuffer16 is  begin    process(Data, En)      begin      if (En = '1') then        Outp <= Data;      else        Outp <= "ZZZZZZZZZZZZZZZZ";      end if;    end process;end behav;
